package Tb;

module mkTb(Empty);
   
   rule hello;
      $display("Hello, world!");
      $finish;
   endrule
   
endmodule

endpackage
